library verilog;
use verilog.vl_types.all;
entity tst_4 is
end tst_4;
