library verilog;
use verilog.vl_types.all;
entity testbench_PC is
end testbench_PC;
