library verilog;
use verilog.vl_types.all;
entity testbench_clock is
end testbench_clock;
