library verilog;
use verilog.vl_types.all;
entity testbench_zero_extend is
end testbench_zero_extend;
