library verilog;
use verilog.vl_types.all;
entity testbench_Adder is
end testbench_Adder;
