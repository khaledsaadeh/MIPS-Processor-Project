library verilog;
use verilog.vl_types.all;
entity tst_5 is
end tst_5;
