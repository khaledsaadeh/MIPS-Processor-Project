library verilog;
use verilog.vl_types.all;
entity tst_6 is
end tst_6;
