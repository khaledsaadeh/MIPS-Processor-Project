library verilog;
use verilog.vl_types.all;
entity testbench_sign_extend is
end testbench_sign_extend;
