library verilog;
use verilog.vl_types.all;
entity testbench_RegisterFile is
end testbench_RegisterFile;
