library verilog;
use verilog.vl_types.all;
entity tst_7 is
end tst_7;
