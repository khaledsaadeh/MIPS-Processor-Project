library verilog;
use verilog.vl_types.all;
entity tst_2 is
end tst_2;
