library verilog;
use verilog.vl_types.all;
entity tst_9 is
end tst_9;
