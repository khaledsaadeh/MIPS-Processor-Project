library verilog;
use verilog.vl_types.all;
entity testbench_Forwarding_unit is
end testbench_Forwarding_unit;
