library verilog;
use verilog.vl_types.all;
entity testbench_control_unit is
end testbench_control_unit;
