library verilog;
use verilog.vl_types.all;
entity Top is
    port(
        PC_VALUE        : in     vl_logic
    );
end Top;
