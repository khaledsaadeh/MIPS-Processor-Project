library verilog;
use verilog.vl_types.all;
entity testbench_mux_2to1 is
end testbench_mux_2to1;
