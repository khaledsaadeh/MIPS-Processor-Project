library verilog;
use verilog.vl_types.all;
entity tst_8 is
end tst_8;
