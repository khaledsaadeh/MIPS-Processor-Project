library verilog;
use verilog.vl_types.all;
entity testbench_IF_ID is
end testbench_IF_ID;
