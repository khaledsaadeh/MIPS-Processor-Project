library verilog;
use verilog.vl_types.all;
entity testbench_shift_left_26bits is
end testbench_shift_left_26bits;
