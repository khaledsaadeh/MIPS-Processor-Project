library verilog;
use verilog.vl_types.all;
entity testbench_memory is
end testbench_memory;
