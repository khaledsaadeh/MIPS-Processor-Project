library verilog;
use verilog.vl_types.all;
entity arethmatic1 is
end arethmatic1;
