library verilog;
use verilog.vl_types.all;
entity tst_1 is
end tst_1;
